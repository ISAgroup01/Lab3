package CONSTANTS is
   constant NumBit : integer := 4;		
end CONSTANTS;
