LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE RISCV_package is
  
  constant nb_i : integer := 32; --Number of bits instruction
  
END PACKAGE;
