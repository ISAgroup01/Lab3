isa01@localhost.localdomain.27352:1612743535