package alu_types is
	type TYPE_OP is (ADD, SUB, BITAND, BITXOR,  FUNCASR);
end alu_types;
